** sch_path: /foss/designs/Workshop_CASS/Módulo_Analógico/Laboratorios/Lab5/Inverter/xschem/inverter.sch
.subckt inverter Vin VDD VSS Vout
*.PININFO Vin:I VDD:B VSS:B Vout:B
M1 Vout Vin VSS VSS nfet_03v3 L=1u W=3u nf=1 m=1
M2 Vout Vin VDD VDD pfet_03v3 L=1u W=3u nf=1 m=1
.ends
