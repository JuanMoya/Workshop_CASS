magic
tech sky130A
timestamp 1761516804
<< nwell >>
rect -153 -9 205 80
rect 95 -10 205 -9
<< nmos >>
rect -85 -160 -70 -110
rect -20 -160 -5 -110
rect 45 -160 60 -110
rect 105 -160 120 -110
<< pmos >>
rect -85 10 -70 60
rect -20 10 -5 60
rect 45 10 60 60
rect 105 10 120 60
<< ndiff >>
rect -135 -127 -85 -110
rect -135 -147 -120 -127
rect -100 -147 -85 -127
rect -135 -160 -85 -147
rect -70 -127 -20 -110
rect -70 -147 -55 -127
rect -35 -147 -20 -127
rect -70 -160 -20 -147
rect -5 -127 45 -110
rect -5 -147 10 -127
rect 30 -147 45 -127
rect -5 -160 45 -147
rect 60 -127 105 -110
rect 60 -147 73 -127
rect 93 -147 105 -127
rect 60 -160 105 -147
rect 120 -127 186 -110
rect 120 -147 135 -127
rect 155 -147 186 -127
rect 120 -160 186 -147
<< pdiff >>
rect -135 43 -85 60
rect -135 23 -120 43
rect -100 23 -85 43
rect -135 10 -85 23
rect -70 43 -20 60
rect -70 23 -55 43
rect -35 23 -20 43
rect -70 10 -20 23
rect -5 43 45 60
rect -5 23 10 43
rect 30 23 45 43
rect -5 10 45 23
rect 60 10 105 60
rect 120 43 185 60
rect 120 23 135 43
rect 155 23 185 43
rect 120 10 185 23
<< ndiffc >>
rect -120 -147 -100 -127
rect -55 -147 -35 -127
rect 10 -147 30 -127
rect 73 -147 93 -127
rect 135 -147 155 -127
<< pdiffc >>
rect -120 23 -100 43
rect -55 23 -35 43
rect 10 23 30 43
rect 135 23 155 43
<< poly >>
rect -85 60 -70 75
rect -20 60 -5 75
rect 45 60 60 76
rect 105 60 120 76
rect -85 -110 -70 10
rect -20 -110 -5 10
rect 45 -110 60 10
rect 105 -110 120 10
rect -85 -175 -70 -160
rect -20 -175 -5 -160
rect 45 -175 60 -160
rect 105 -175 120 -160
<< locali >>
rect -136 94 220 114
rect -125 43 -95 51
rect -125 23 -120 43
rect -100 23 -95 43
rect -125 15 -95 23
rect -60 43 -30 51
rect 10 50 30 94
rect -60 23 -55 43
rect -35 23 -30 43
rect -60 15 -30 23
rect 5 43 35 50
rect 5 23 10 43
rect 30 23 35 43
rect 5 15 35 23
rect 130 43 160 51
rect 130 23 135 43
rect 155 23 160 43
rect 130 15 160 23
rect -120 -40 -100 15
rect -55 -3 -35 15
rect 135 -3 155 15
rect -55 -20 155 -3
rect 200 -40 231 -28
rect -120 -57 231 -40
rect -55 -118 -36 -57
rect 200 -66 231 -57
rect 10 -97 155 -75
rect 10 -118 30 -97
rect 135 -118 155 -97
rect -125 -127 -95 -118
rect -125 -147 -120 -127
rect -100 -147 -95 -127
rect -125 -155 -95 -147
rect -60 -127 -30 -118
rect -60 -147 -55 -127
rect -35 -147 -30 -127
rect -60 -155 -30 -147
rect 5 -127 35 -118
rect 5 -147 10 -127
rect 30 -147 35 -127
rect 5 -155 35 -147
rect 68 -127 98 -118
rect 68 -147 73 -127
rect 93 -147 98 -127
rect 68 -155 98 -147
rect 130 -127 160 -118
rect 130 -147 135 -127
rect 155 -147 160 -127
rect 130 -155 160 -147
rect -120 -185 -99 -155
rect 73 -185 94 -155
rect -135 -205 220 -185
<< labels >>
rlabel poly -85 -175 -70 -160 5 A
port 1 s
rlabel poly -20 -175 -5 -160 5 B
port 2 s
rlabel poly 45 -175 60 -160 5 C
port 3 s
rlabel poly 105 -175 120 -160 5 D
port 4 s
rlabel locali 200 -66 231 -28 3 Q
port 5 e
rlabel locali -136 94 220 114 7 VPWR
port 6 w
rlabel locali -135 -205 220 -185 7 VGND
port 7 w
<< end >>
