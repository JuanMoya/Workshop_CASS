** sch_path: /foss/designs/Workshop_CASS/Modulo_Analogico/Laboratorios/Lab2/inv_tb.sch
**.subckt inv_tb
x1 Vin VDD VSS Vout inverter
C1 Vout VSS 100f m=1
V1 VSS GND 0
V2 VDD VSS 3.3
Vin Vin VSS PULSE(0 3.3 0 5n 5n 1u 2u)
**** begin user architecture code

.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/smbb000149.ngspice typical



*Parameters

.options TEMP = 27

.control
*Transient analysis
tran 0.1n 10u
save all
let VP=3.3
let per10 = Vp*0.1
let per50 = Vp*0.5
let per90 = Vp*0.9
meas tran t_rise  TRIG v(Vout) VAL=per10 rise=2  TARG v(Vout) VAL=per90 rise=2
meas tran t_fall  TRIG v(Vout) VAL=per90 fall=2  TARG v(Vout) VAL=per10 fall=2
meas tran t_delay  TRIG v(Vin) VAL=per50 rise=1 TARG v(Vout) VAL=per50 fall=1
echo tran measurements
print t_delay
print t_rise
print t_fall
echo

set filetype=ascii
write results.txt v(Vin) v(Vout) time
.endc
.end


**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /foss/designs/Workshop_CASS/Modulo_Analogico/Laboratorios/Lab2/inverter.sym
** sch_path: /foss/designs/Workshop_CASS/Modulo_Analogico/Laboratorios/Lab2/inverter.sch
.subckt inverter Vin VDD VSS Vout
*.ipin Vin
*.iopin VDD
*.iopin VSS
*.iopin Vout
XM1 Vout Vin VSS VSS nfet_03v3 L=1u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 Vout Vin VDD VDD pfet_03v3 L=1u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
