** sch_path: /foss/designs/Workshop_CASS/Modulo_Analogico/Laboratorios/Lab4/current_mirror_improved.sch
**.subckt current_mirror_improved
Vdd v_dd GND 3.3
Ibias v_dd v_gs 20u
Vout1 out1 GND 0.6
Vout2 out2 GND 0.6
Vout3 out3 GND 0.6
.save v(out1)
.save v(out2)
.save v(out3)
.save v(v_gs)
Viout1 out1 net1 0
.save i(viout1)
Viout2 out2 net2 0
.save i(viout2)
Viout3 out3 net3 0
.save i(viout3)
XM1 v_gs v_gs GND GND nfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 net1 v_gs GND GND nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 net2 v_gs GND GND nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net3 v_gs GND GND nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
**** begin user architecture code


.temp 27
.control
save all

op
write current_mirror_improved.raw
dc Vout1 0 3.3 10m
plot i(viout1) vs v(out1)
dc Vout2 0 3.3 10m
plot i(viout2) vs v(out2)
dc Vout3 0 3.3 10m
plot i(viout3) vs v(out3)

.endc



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/smbb000149.ngspice typical

**** end user architecture code
**.ends
.GLOBAL GND
.end
