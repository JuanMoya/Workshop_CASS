* NGSPICE file created from 3_stage_RO.ext - technology: gf180mcuD

.subckt 3_stage_RO VDD VSS n1
X0 a_1240_314# a_240_314# VDD.t3 VDD.t2 pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=1u
X1 a_1240_314# a_240_314# VSS.t1 VSS.t0 nfet_03v3 ad=1.83p pd=7.22u as=1.83p ps=7.22u w=3u l=1u
X2 a_240_314# n1.t2 VDD.t1 VDD.t0 pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=1u
X3 a_240_314# n1.t3 VSS.t5 VSS.t4 nfet_03v3 ad=1.83p pd=7.22u as=1.83p ps=7.22u w=3u l=1u
X4 n1.t0 a_1240_314# VSS.t3 VSS.t2 nfet_03v3 ad=1.83p pd=7.22u as=1.83p ps=7.22u w=3u l=1u
X5 n1.t1 a_1240_314# VDD.t5 VDD.t4 pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=1u
R0 VDD.t2 VDD.n2 764.841
R1 VDD.t0 VDD.n4 764.841
R2 VDD.n5 VDD.t0 379.233
R3 VDD.n2 VDD.t4 376.712
R4 VDD.n4 VDD.t2 376.712
R5 VDD.n1 VDD.n0 3.12818
R6 VDD VDD.n5 2.94908
R7 VDD.n3 VDD.n0 2.67312
R8 VDD.n2 VDD.n1 2.5205
R9 VDD.n4 VDD.n3 2.5205
R10 VDD.n3 VDD.t3 2.0205
R11 VDD.n1 VDD.t5 2.0205
R12 VDD.n5 VDD.t1 2.0205
R13 VDD VDD.n0 0.178839
R14 VSS.t0 VSS.n2 1250.57
R15 VSS.t4 VSS.n4 1250.57
R16 VSS.n5 VSS.t4 596.008
R17 VSS.n2 VSS.t2 593.928
R18 VSS.n4 VSS.t0 593.928
R19 VSS.n1 VSS.n0 3.12779
R20 VSS VSS.n5 2.96854
R21 VSS.n3 VSS.n0 2.67272
R22 VSS.n3 VSS.t1 2.1005
R23 VSS.n1 VSS.t3 2.1005
R24 VSS.n5 VSS.t5 2.1005
R25 VSS.n2 VSS.n1 2.0805
R26 VSS.n4 VSS.n3 2.0805
R27 VSS VSS.n0 0.159748
R28 n1.n0 n1.t2 27.7092
R29 n1.n0 n1.t3 27.157
R30 n1.n2 n1.n0 6.4625
R31 n1.n2 n1.n1 4.5005
R32 n1.n1 n1.t1 3.98765
R33 n1.n1 n1.t0 3.70386
R34 n1 n1.n2 0.0059
C0 a_240_314# VDD 0.92277f
C1 a_1240_314# VDD 0.91181f
C2 n1 VDD 0.68039f
C3 a_1240_314# a_240_314# 0.4723f
C4 n1 a_240_314# 0.87652f
C5 n1 a_1240_314# 0.87363f
C6 n1 VSS 2.47638f
C7 VDD VSS 8.71481f
C8 a_1240_314# VSS 1.60183f
C9 a_240_314# VSS 1.59372f
.ends

