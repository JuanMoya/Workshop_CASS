** sch_path: /foss/designs/Workshop_CASS/Módulo_Analógico/Laboratorios/Lab5/Inverter/pex/inverter_tb_none.sch
**.subckt inverter_tb_none
C1 Vout VSS 1f m=1
V1 VSS GND 0
V2 VDD VSS 3.3
Vin Vin VSS 0
X1 Vin VDD VSS Vout inverter
**** begin user architecture code

.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/smbb000149.ngspice typical



.include /foss/designs/Workshop_CASS/Módulo_Analógico/Laboratorios/Lab5/Inverter/pex/inverter.spice
.control
dc Vin 0 3.3 0.01
plot v(Vout)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
